`timescale 1ns / 1ps
module IM_unit(
    input [7:0] Addr,		//ָ��洢����ַ���� 
    output [31:0]  instruction// �Ĵ�����ֵ
);
    reg [31:0] IM [0:255]; // �Ĵ�����
    assign instruction=IM[Addr];
    integer i;
    initial begin
        IM[0]<=32'h00000000;    //0000
        IM[1]<=32'h24010008;    //0004
        IM[2]<=32'h34020002;    //0008
        IM[3]<=32'h00411820;    //000c
        IM[4]<=32'h00622822;    //0010
        IM[5]<=32'h00a22024;    //0014
        IM[6]<=32'h00824025;    //0018
        IM[7]<=32'h00084040;    //001c
        IM[8]<=32'h1501fffe;    //0020
        IM[9]<=32'h28460004;    //0024
        IM[10]<=32'h28c7ffff;   //0028
        IM[11]<=32'h2cc6ffff;   //002c
        IM[12]<=32'h20e70008;   //0030
        IM[13]<=32'h10e1fffe;   //0034
        IM[14]<=32'h2001ffff;   //0038
        IM[15]<=32'h254a0001;   //003c
        IM[16]<=32'h0540fffe;   //0040
        IM[17]<=32'h304b0002;   //0044
        IM[18]<=32'h0c000038;   //0048 jal
        IM[19]<=32'h004b4026;   //004c
        IM[20]<=32'h00cb4027;   //0050
        IM[21]<=32'h010b4021;   //0054
        IM[22]<=32'h01064023;   //0058
        IM[23]<=32'h00010842;   //005c
        IM[24]<=32'h00084083;   //0060
        IM[25]<=32'h3c090007;   //0064
        IM[26]<=32'h0028502a;   //0068
        IM[27]<=32'h0028502b;   //006c
        IM[28]<=32'h00c82004;   //0070
        IM[29]<=32'h20840001;   //0074
        IM[30]<=32'h1880fffe;   //0078
        IM[31]<=32'h05100017;   //007c
        IM[32]<=32'h2042ffff;   //0080
        IM[33]<=32'h1c40fffe;   //0084
        IM[34]<=32'h216bffff;   //0088
        IM[35]<=32'h0561fffe;   //008c
        IM[36]<=32'h04110012;   //0090
        IM[37]<=32'h00e86006;   //0094
        IM[38]<=32'h00e86007;   //0098
        IM[39]<=32'h71801021;   //009c
        IM[40]<=32'h000c6100;   //00a0
        IM[41]<=32'h71801021;   //00a4
        IM[42]<=32'h71001020;   //00a8
        IM[43]<=32'h000841c2;   //00ac
        IM[44]<=32'h71001020;   //00b0
        IM[45]<=32'h70430802;   //00b4
        IM[46]<=32'h004b0018;   //00b8
        IM[47]<=32'h004b0019;   //00bc
        IM[48]<=32'h00e5001a;   //00c0
        IM[49]<=32'h0027001b;   //00c4
        IM[50]<=32'h00002010;   //00c8
        IM[51]<=32'h00003012;   //00cc
        IM[52]<=32'h00a00011;   //00d0
        IM[53]<=32'h00200013;   //00d4
        IM[54]<=32'h0800003a;   //00d8
        IM[55]<=32'h03e00008;   //00dc
        IM[56]<=32'h23fe0000;   //00e0 addi
        IM[57]<=32'h03c0f809;   //00e4 jalr
        IM[58]<=32'h714b0000;   //00e8
        IM[59]<=32'h714b0001;   //00ec
        IM[60]<=32'h70a60004;   //00f0
        IM[61]<=32'h714b0005;   //00f4
        IM[62]<=32'haca80000;   //00f8
        IM[63]<=32'ha4a80004;   //00fc
        IM[64]<=32'ha0a80008;   //0100
        IM[65]<=32'h8ca10000;   //0104
        IM[66]<=32'h20210000;   //0108
        IM[67]<=32'h8ca10004;   //010c
        IM[68]<=32'h20210000;   //0110
        IM[69]<=32'h8ca10008;   //0114
        IM[70]<=32'h20210000;   //0118
        IM[71]<=32'h84a10000;   //011c
        IM[72]<=32'h20210000;   //0120
        IM[73]<=32'h94a10000;   //0124
        IM[74]<=32'h20210000;   //0128
        IM[75]<=32'h80a10000;   //012c
        IM[76]<=32'h20210000;   //0130
        IM[77]<=32'h90a10000;   //0134
        IM[78]<=32'h20210000;   //0138
        IM[79]<=32'h3981ffff;   //013c
        //IM[80]<=32'h;
        //IM[81]<=32'h;
        for(i=80;i<256;i=i+1)
            IM[i]<=0;
    end
endmodule 
